
`include "apb_top.sv"
`include "apb_test.sv"


module apb_testbench_top;

  bit PCLK;                //clock signal declaration
  bit RESET;                //reset signal declaration

  //interface instance
   apb_intf intf (PCLK,RESET);
  //   apb_intf intf (PCLK,RESET,sysbus,PRDATA);
  //DUT instance, interface signals are connected to the DUT ports
  top_apb DUT (
    .PCLK(intf.PCLK),
    .RESET(intf.RESET),
    .sysbus(intf.sysbus),
    .PRDATA(intf.RDATA)
   );

  always #5 PCLK = ~PCLK;   //clock generation
  //reset Generation
  initial begin
    RESET = 1;
    #5 RESET =0;
  end

  //passing the interface handle to lower heirarchy using set method and enabling the wave dump
  initial begin 
    uvm_config_db#(virtual apb_intf)::set(uvm_root::get(),"*","intf",intf);
    //enable wave dump
    $dumpfile("dump.vcd"); 
    $dumpvars;
  end
  
  initial begin 
    run_test();
  end
  
endmodule