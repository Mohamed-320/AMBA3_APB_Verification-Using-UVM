
/*************** Simple Bridge/Slave DUT***************/
module top_apb(PCLK,RESET,sysbus,PRDATA);
input PCLK,RESET;
input [20:0] sysbus;
output reg [7:0] PRDATA;
wire PSEL,PENABLE,PWRITE;
wire [7:0] PADDR;
wire [7:0] PWDATA;

apb_bridge DUT1( .PCLK(PCLK),
                 .RESET(RESET),
                 .PENABLE(PENABLE), 
                 .PSEL(PSEL), 
                 .PWRITE(PWRITE), 
                 .PADDR(PADDR),
                 .PWDATA(PWDATA), 
                 .PRDATA(PRDATA),
                 .system_bus(sysbus));

apb_slave DUT2( .PCLK(PCLK),
                .RESET(RESET),
                .PENABLE(PENABLE), 
                .PSEL(PSEL), 
                .PWRITE(PWRITE),
                .PADDR(PADDR), 
                .PWDATA(PWDATA), 
                .PRDATA(PRDATA));
endmodule
