

/***************Monitor samples the DUT signals through the virtual interface and converts the signal level activity to the transaction level**************/
`ifndef APB_MONITOR
`define APB_MONITOR

import uvm_pkg::*;        // Standard UVM pkg
`include "uvm_macros.svh" //Standard UVM macros
`include "apb_driver.sv"

class apb_monitor extends uvm_monitor;

virtual apb_intf intf;  // virtual interface
uvm_analysis_port#(apb_seq_item) item_collected_port; //analysis port
apb_seq_item trans_collected; //seq_item handle, used as a place holder for sampled signal activity (to capture transaction info)

    `uvm_component_utils(apb_monitor)

      function new(string name,uvm_component parent);
         super.new(name,parent);
         trans_collected=new();
         item_collected_port=new("item_collected_port",this);
      endfunction : new

       function void build_phase(uvm_phase phase);
         super.build_phase(phase);
         if(!uvm_config_db#(virtual apb_intf)::get(this,"","intf",intf))`uvm_fatal("No interface",{"virtual interface must be set for: ",get_full_name(),".intf"});
       endfunction : build_phase

  virtual task run_phase(uvm_phase phase);
  forever begin
   @(posedge intf.MONITOR.PCLK);
   trans_collected.sysbus=intf.monitor_cb.sysbus;

   @(posedge intf.MONITOR.PCLK);
   trans_collected.PRDATA=intf.monitor_cb.PRDATA;

   item_collected_port.write(trans_collected);
   end
  endtask: run_phase
endclass : apb_monitor

`endif