
/************************** The test defines the test scenario for the testbench **********************************/  
`ifndef APB_TEST
`define APB_TEST

import uvm_pkg::*;        // Standard UVM pkg
`include "uvm_macros.svh" //Standard UVM macros
`include "apb_env.sv"

class apb_test extends uvm_test;
apb_env env;

`uvm_component_utils(apb_test)
 function new(string name="apb_test",uvm_component parent=null);
  super.new(name,parent);
 endfunction : new

 virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    // Create the env
    env = apb_env::type_id::create("env", this);
  endfunction : build_phase

  task run_phase(uvm_phase phase);
      phase.raise_objection(this);
      seq.start(env.agent.sequencer);
      phase.drop_objection(this);
  endtask : run_phase
endclass 
`endif